module and_gate
    (
        input logic A,
        input logic B,
        input logic C,
    );

    assign Y = A & B;

endmodule
